
module Nand2Tetris
(
	input         clk,
	input         reset,

	// input         pal,
	input         scandouble,

	output reg    ce_pix,

	output reg    HBlank,
	output reg    HSync,
	output reg    VBlank,
	output reg    VSync,

	output  [7:0] video
);



endmodule
